`timescale 1ns / 1ps
// <111550168>

/** [Prerequisite] pipelined (Lab 3), forwarding, hazard_detection
 * This module is the pipelined MIPS processor "similar to" FIGURE 4.60 (control hazard is not solved).
 * You can implement it by any style you want, as long as it passes testbench.
 */

module pipelined #(
    parameter integer TEXT_BYTES = 1024,        // size in bytes of instruction memory
    parameter integer TEXT_START = 'h00400000,  // start address of instruction memory
    parameter integer DATA_BYTES = 1024,        // size in bytes of data memory
    parameter integer DATA_START = 'h10008000   // start address of data memory
) (
    input clk,  // clock
    input rstn  // negative reset
);

    /** [step 0] Copy from Lab 3

    /* Instruction Memory */
    wire [31:0] instr_mem_address, instr_mem_instr;
    instr_mem #(
        .BYTES(TEXT_BYTES),
        .START(TEXT_START)
    ) instr_mem (
        .address(instr_mem_address),
        .instr  (instr_mem_instr)
    );

    /* Register Rile */
    wire [4:0] reg_file_read_reg_1, reg_file_read_reg_2, reg_file_write_reg;
    wire reg_file_reg_write;
    wire [31:0] reg_file_write_data, reg_file_read_data_1, reg_file_read_data_2;
    reg_file reg_file (
        .clk        (~clk),                  // only write when negative edge
        .rstn       (rstn),
        .read_reg_1 (reg_file_read_reg_1),
        .read_reg_2 (reg_file_read_reg_2),
        .reg_write  (reg_file_reg_write),
        .write_reg  (reg_file_write_reg),
        .write_data (reg_file_write_data),
        .read_data_1(reg_file_read_data_1),//output
        .read_data_2(reg_file_read_data_2)//output
    );

    /* ALU */
    wire [31:0] alu_a, alu_b, alu_result;
    wire [3:0] alu_ALU_ctl;
    wire alu_zero, alu_overflow;
    alu alu (
        .a       (alu_a),
        .b       (alu_b),
        .ALU_ctl (alu_ALU_ctl),
        .result  (alu_result),
        .zero    (alu_zero),
        .overflow(alu_overflow)
    );
    //assign alu_a = ID_EX_read_data_1;
    //assign alu_b = (ID_EX_alu_src) ? ID_EX_sign_extend : ID_EX_read_data_2;
    assign alu_ALU_ctl = alu_control_operation;

    /* Data Memory */
    wire data_mem_mem_read, data_mem_mem_write;
    wire [31:0] data_mem_address, data_mem_write_data, data_mem_read_data;
    data_mem #(
        .BYTES(DATA_BYTES),
        .START(DATA_START)
    ) data_mem (
        .clk       (~clk),                 // only write when negative edge
        .mem_read  (data_mem_mem_read),
        .mem_write (data_mem_mem_write),
        .address   (data_mem_address),
        .write_data(data_mem_write_data),
        .read_data (data_mem_read_data) //output
    );
    assign data_mem_mem_read = EX_MEM_mem_read;
    assign data_mem_mem_write = EX_MEM_mem_write;
    assign data_mem_address = EX_MEM_alu_result;
    assign data_mem_write_data = EX_MEM_read_data_2;
    

    /* ALU Control */
    wire [1:0] alu_control_alu_op;
    wire [5:0] alu_control_funct;
    wire [3:0] alu_control_operation;
    alu_control alu_control (
        .alu_op   (alu_control_alu_op),
        .funct    (alu_control_funct),
        .operation(alu_control_operation)
    );
    assign alu_control_alu_op = ID_EX_alu_op;
    assign alu_control_funct = ID_EX_sign_extend[5:0];

    /* (Main) Control */
    wire [5:0] control_opcode;
    wire [5:0] control_funct;
    // Execution/address calculation stage control lines
    wire control_reg_dst, control_alu_src;
    wire [1:0] control_alu_op;
    // Memory access stage control lines
    wire control_branch, control_mem_read, control_mem_write;
    // Wire-back stage control lines
    wire control_reg_write, control_mem_to_reg;
    control control (
        .opcode    (control_opcode),//input
        .funct     (control_funct),//input
        //.stall     (stall),//input
        .reg_dst   (control_reg_dst),
        .alu_src   (control_alu_src),
        .mem_to_reg(control_mem_to_reg),
        .reg_write (control_reg_write),
        .mem_read  (control_mem_read),
        .mem_write (control_mem_write),
        .branch    (control_branch),
        .alu_op    (control_alu_op)
    );

    /** [step 1] Instruction fetch (IF)
     * 1. We need a register to store PC (acts like pipeline register).
     * 2. Wire pc to instruction memory.
     * 3. Implement an adder to calculate PC+4. (combinational)
     *    Hint: use "+" operator.
     * 4. Update IF/ID pipeline registers, and reset them @(negedge rstn)
     *    a. fetched instruction
     *    b. PC+4
     *    Hint: What else should be done when reset?
     *    Hint: Update of PC can be handle later in MEM stage.
     */
    // 1.
    reg [31:0] pc;  // DO NOT change this line
    // 2.
    assign instr_mem_address = pc;
    // 3.
    wire [31:0] pc_4;
    assign pc_4 = pc +4;
    // 4.
    reg [31:0] IF_ID_instr, IF_ID_pc_4;
    always @(posedge clk)
        if (rstn && IF_ID_write) begin //rstn is 1 means it's safe to update new value to register
            IF_ID_instr <=  instr_mem_instr;  // a.
            IF_ID_pc_4  <= pc_4;  // b.
        end
    always @(negedge rstn) begin
        IF_ID_instr <= 0;  // a.
        IF_ID_pc_4  <= 0;  // b.
    end


    /** [step 2] Instruction decode and register file read (ID)
     * From top to down in FIGURE 4.51: (instr. refers to the instruction from IF/ID)
     * 1. Generate control signals of the instr. (as Lab 2)
     * 2. Read desired registers (from register file) in the instr.
     * 3. Calculate sign-extended immediate from the instr.
     * 4. Update ID/EX pipeline registers, and reset them @(negedge rstn)
     *    a. Control signals (WB, MEM, EX)
     *    b. ??? (something from IF/ID)
     *    c. Data read from register file
     *    d. Sign-extended immediate
     *    e. ??? & ??? (WB stage needs to know which reg to write)
     */
    assign control_opcode = IF_ID_instr[31:26];
    assign control_funct = IF_ID_instr[5:0];
    assign reg_file_read_reg_1= IF_ID_instr[25:21];
    assign reg_file_read_reg_2 = IF_ID_instr[20:16];
    // 3.
    wire[31:0] sign_extend;
    assign sign_extend = {{16{IF_ID_instr[15]}}, IF_ID_instr[15:0]};

    //ID stage  setup
    reg [31:0] ID_EX_sign_extend;
    reg [4:0] ID_EX_rs, ID_EX_rt, ID_EX_rd;
    reg ID_EX_reg_write,ID_EX_mem_to_reg; //WB
    reg ID_EX_mem_read, ID_EX_mem_write;
    //reg ID_EX_branch; //M
    reg ID_EX_alu_src, ID_EX_reg_dst; //EX
    reg [1:0] ID_EX_alu_op; //EX
    reg [31:0] ID_EX_read_data_1, ID_EX_read_data_2;
    reg [31:0]ID_EX_pc_4;


    always @(posedge clk or negedge rstn) begin
        if (!rstn) begin
            // Reset ID/EX pipeline registers
            ID_EX_sign_extend <= 0;
            ID_EX_rs <= 0;
            ID_EX_rt <= 0;
            ID_EX_rd <= 0;
            ID_EX_reg_write <= 0;
            ID_EX_mem_to_reg <= 0;
            ID_EX_mem_read <= 0;
            ID_EX_mem_write <= 0;
            //ID_EX_branch <= 0;
            ID_EX_alu_src <= 0;
            ID_EX_reg_dst <= 0;
            ID_EX_alu_op <= 0;
            ID_EX_read_data_1 <= 0;
            ID_EX_read_data_2 <= 0;
            ID_EX_pc_4 <= 0;
        end else begin
            // Pass decoded data to EX stage
            ID_EX_sign_extend <=sign_extend;
            ID_EX_rs <= reg_file_read_reg_1;
            ID_EX_rt <= IF_ID_instr[20:16]; //TODO: R-fromat or I-format
            ID_EX_rd <= IF_ID_instr[15:11];  // destination register
            ID_EX_reg_write <= stall? 0:control_reg_write;
            ID_EX_mem_to_reg <= stall? 0:control_mem_to_reg;
            ID_EX_mem_read <= stall? 0:control_mem_read;
            ID_EX_mem_write <= stall? 0:control_mem_write;
            //ID_EX_branch <= control_branch;
            ID_EX_alu_src <= stall? 0:control_alu_src;
            ID_EX_reg_dst <= stall? 0:control_reg_dst;
            ID_EX_alu_op <= control_alu_op;
            ID_EX_read_data_1 <= reg_file_read_data_1;
            ID_EX_read_data_2 <= reg_file_read_data_2;
            ID_EX_pc_4 <= IF_ID_pc_4;
        end
    end

    always @(posedge clk)
        if (rstn) begin
        pc <=  ID_branch_taken? ID_branch_target :(pc_write? pc_4:pc);
        end
    always @(negedge rstn) begin
        pc <= 32'h00400000;
    end

    /** [step 3] Execute or address calculation (EX)
     * From top to down in FIGURE 4.51
     * 1. Calculate branch target address from sign-extended immediate.
     * 2. Select correct operands of ALU like in Lab 2.
     * 3. Wire control signals to ALU control & ALU like in Lab 2.
     * 4. Select correct register to write.
     * 5. Update EX/MEM pipeline registers, and reset them @(negedge rstn)
     *    a. Control signals (WB, MEM)
     *    b. Branch target address
     *    c. ??? (What information dose MEM stage need to determine whether to branch?)
     *    d. ALU result
     *    e. ??? (What information does MEM stage need when executing Store?)
     *    f. ??? (WB stage needs to know which reg to write)
     */

    //  EX Stage
    reg [31:0] EX_MEM_alu_result;
    //reg EX_MEM_branch_target;
    reg EX_MEM_zero_flag;
    reg EX_MEM_reg_write, EX_MEM_mem_to_reg; // WB
    reg EX_MEM_mem_read, EX_MEM_mem_write;
    //reg EX_MEM_branch; // MEM
    reg [4:0] EX_MEM_write_reg;
    reg [31:0] EX_MEM_read_data_2;
    reg [31:0]EX_MEM_pc_4;


    always @(posedge clk or negedge rstn) begin
        if (!rstn) begin
            EX_MEM_alu_result <= 0;
            //EX_MEM_branch_target <= 0;
            EX_MEM_zero_flag <= 0;
            EX_MEM_reg_write <= 0;
            EX_MEM_mem_read <= 0;
            EX_MEM_mem_write <= 0;
            //EX_MEM_branch <= 0;
            EX_MEM_mem_to_reg <= 0;
            EX_MEM_write_reg <= 0;
            EX_MEM_read_data_2 <= 0;
            EX_MEM_pc_4 <= 0;
        end else begin
            // Calculate ALU result, branch target, etc.
            EX_MEM_alu_result <= alu_result;  //
            //EX_MEM_branch_target <= ID_EX_pc_4 + (ID_EX_sign_extend << 2);  // Branch target 
            EX_MEM_zero_flag <= alu_zero;
            EX_MEM_reg_write <= ID_EX_reg_write;
            EX_MEM_mem_read <= ID_EX_mem_read;
            EX_MEM_mem_write <= ID_EX_mem_write;
            //EX_MEM_branch <= ID_EX_branch;
            EX_MEM_mem_to_reg <= ID_EX_mem_to_reg;
            EX_MEM_write_reg <= write_reg_address;  // Choose register to write
            EX_MEM_read_data_2 <= ID_EX_read_data_2;
            EX_MEM_pc_4 <= ID_EX_pc_4;
        end
    end
    wire [31:0]write_reg_address;
    assign write_reg_address = ID_EX_reg_dst ? ID_EX_rd : ID_EX_rt;



    /** [step 4] Memory access (MEM)
     * From top to down in FIGURE 4.51
     * 1. Decide whether to branch or not.
     * 2. Wire address & data to write
     * 3. Wire control signal of read/write
     * 4. Update MEM/WB pipeline registers, and reset them @(negedge rstn)
     *    a. Control signals (WB)
     *    b. ???
     *    c. ???
     *    d. ???
     * 5. Update PC.
     */
    //wire pc_src;
    //assign pc_src = EX_MEM_branch && EX_MEM_zero_flag; 

    // Memory Access (MEM) Stage
    reg [31:0] MEM_WB_write_data, MEM_WB_address;
    reg MEM_WB_reg_write, MEM_WB_mem_to_reg;
    reg [4:0] MEM_WB_write_reg;

    always @(posedge clk or negedge rstn) begin
        if (!rstn) begin
            MEM_WB_write_data <= 0;
            MEM_WB_address <= 0;
            MEM_WB_reg_write <= 0;
            MEM_WB_mem_to_reg <= 0;
            MEM_WB_write_reg <= 0;
            pc <= 32'h00400000;
        end 
        else begin
            // Decide whether to branch
            //pc <= pc_write? pc_4: (pc_src? EX_MEM_branch_target :pc);  // change to ID stage

            // Data memory operations
            MEM_WB_write_data <= data_mem_read_data;  // Data from memory
            MEM_WB_address <= EX_MEM_alu_result;
            MEM_WB_reg_write <= EX_MEM_reg_write;
            MEM_WB_mem_to_reg <= EX_MEM_mem_to_reg;
            MEM_WB_write_reg <= EX_MEM_write_reg;
        end
    end


    /** [step 5] Write-back (WB)
     * From top to down in FIGURE 4.51
     * 1. Wire RegWrite of register file.
     * 2. Select the data to write into register file.
     * 3. Select which register to write.
     */

    assign reg_file_reg_write = MEM_WB_reg_write;//enable
    assign reg_file_write_data = MEM_WB_mem_to_reg ? MEM_WB_write_data : MEM_WB_address; //lwsw:r-format,i-format
    assign reg_file_write_reg = MEM_WB_write_reg;
    


    //lab4
    /** [step 2] Connect Forwarding unit
     * 1. add `ID_EX_rs` into ID/EX stage registers
     * 2. Use a mux to select correct ALU operands according to forward_A/B
     *    Hint don't forget that alu_b might be sign-extended immediate!
     */
    wire [1:0] forward_A, forward_B;
    forwarding forwarding (
        .ID_EX_rs        (ID_EX_rs),
        .ID_EX_rt        (ID_EX_rt),
        .EX_MEM_reg_write(EX_MEM_reg_write),
        .EX_MEM_rd       (EX_MEM_write_reg),//
        .MEM_WB_reg_write(MEM_WB_reg_write),
        .MEM_WB_rd       (MEM_WB_write_reg),//
        .forward_A       (forward_A),
        .forward_B       (forward_B)
    );

    assign alu_a = (forward_A == 2'b01) ? reg_file_write_data : //328
                   (forward_A == 2'b10) ? EX_MEM_alu_result  : ID_EX_read_data_1;

    assign alu_b = (forward_B == 2'b01) ? reg_file_write_data :
                    (forward_B == 2'b10) ? EX_MEM_alu_result  :
                    (ID_EX_alu_src) ? ID_EX_sign_extend :ID_EX_read_data_2; //TODO

    /** [step 4] Connect Hazard Detection unit
     * 1. use `pc_write` when updating PC
     * 2. use `IF_ID_write` when updating IF/ID stage registers
     * 3. use `stall` when updating ID/EX stage registers
     */
    wire cur_branch, pre_load, pre_r_format;
    hazard_detection hazard_detection (
        .ID_EX_mem_read(ID_EX_mem_read),
        .ID_EX_rd      (write_reg_address),
        .IF_ID_rs      (IF_ID_instr[25:21]),
        .IF_ID_rt      (IF_ID_instr[20:16]),
        .cur_branch    (cur_branch),
        //.EX_MEM_alu_result(EX_MEM_alu_result),
        .EX_MEM_mem_read(EX_MEM_mem_read),
        //.pre_r_format  (pre_r_format),
        //.pre_load      (pre_load),  
        .pc_write      (pc_write),            // implicitly declared
        .IF_ID_write   (IF_ID_write),         // implicitly declared
        .stall         (stall)                // implicitly declared
    );

    //assign pre_r_format = (IF_ID_instr == 6'b000000);//TODO
    //assign pre_load = (IF_ID_instr == 6'b100011);
    assign cur_branch = (IF_ID_instr[31:26] == 6'b000100); // beq instruction

    /** [step 5] Control Hazard
     * This is the most difficult part since the textbook does not provide enough information.
     * By reading p.377-379 "Reducing the Delay of Branches",
     * we can disassemble this into the following steps:
     * 1. Move branch target address calculation & taken or not from EX to ID
     * 2. Move branch decision from MEM to ID//
     * 3. Add forwarding for registers used in branch decision from EX/MEM
     * 4. Add stalling:
          branch read registers right after an ALU instruction writes it -> 1 stall
          branch read registers right after a load instruction writes it -> 2 stalls
     */
     //??�判?��branch??��?��??�instruction?��?��?��r-format??�是lw => hazard_detection
     // Branch target address calculation in ID stage
    wire [31:0] ID_branch_target;
    assign ID_branch_target = IF_ID_pc_4 + (sign_extend << 2);

    wire [31:0]branch_a, branch_b;
    assign branch_a = (branch_forward_A == 2'b10)?  EX_MEM_alu_result:
                      (branch_forward_A == 2'b01)?  reg_file_write_data : reg_file_read_data_1;
    assign branch_b = (branch_forward_B == 2'b10)?  EX_MEM_alu_result:
                      (branch_forward_B == 2'b01)?  reg_file_write_data : reg_file_read_data_2;
    // Branch decision in ID stage
    wire ID_branch_taken;
    assign ID_branch_taken = (IF_ID_instr[31:26]==6'b000100) && (branch_a == branch_b);//要�?�麼?��??�branch??�第�??��?��?�第二�?��?�是?��來自mem??��?�是exe??��?��?��?�forwarding，�?�是forwarding?��?��ex stage�?
    
    wire[1:0] branch_forward_A, branch_forward_B;
    branch_forwarding branch_forwarding (
    .IF_ID_rs        (IF_ID_instr[25:21]),          // inputs are pipeline registers relate to forwarding
    .IF_ID_rt        (IF_ID_instr[20:16]),
    .EX_MEM_reg_write(EX_MEM_reg_write),
    .EX_MEM_rd       (EX_MEM_write_reg),
    .MEM_WB_reg_write(MEM_WB_reg_write),
    .MEM_WB_rd       (MEM_WB_write_reg),
    .cur_branch      (cur_branch),
    //.pre_r_format    (pre_r_format),
    .branch_forward_A   (branch_forward_A),         // ALU operand is from: 00:ID/EX, 10: EX/MEM, 01:MEM/WB
    .branch_forward_B   (branch_forward_B)
    );

    //sw_forwarding sw_forwarding (
    //.EX_MEM_rs        (EX_MEM_alu_result),          // inputs are pipeline registers relate to forwarding
    //.EX_MEM_rt        (EX_MEM_write_reg),
    //.MEM_WB_reg_write(MEM_WB_reg_write),
    //.MEM_WB_rd       (MEM_WB_write_reg), //MEM_WB_write_reg?
    //.sw_forward_A       (sw_forward_A),         // ALU operand is from: 00:ID/EX, 10: EX/MEM, 01:MEM/WB
    //.sw_forward_B       (sw_forward_B)
    //);


endmodule  // pipelined
